module test;

endmodule
