module test;
sss
endmodule
